module sevenseg(
input [3:0] data,
input blank,
input minus, 
output reg [7:0] HEX
);

always @(blank, minus, data[3:0])
casex ({blank, minus, data[3:0]})
  6'b1xxxxx: HEX[7:0] = 8'b11111111;     // blank
  6'b01xxxx: HEX[7:0] = 8'b10111111;     // minus
  6'b001111: HEX[7:0] = 8'b10001110;     // F
  6'b001110: HEX[7:0] = 8'b10000110;     // E
  6'b001101: HEX[7:0] = 8'b10100001;     // D
  6'b001100: HEX[7:0] = 8'b11000110;     // C
  6'b001011: HEX[7:0] = 8'b10000011;     // B
  6'b001010: HEX[7:0] = 8'b10001000;     // A
  6'b001001: HEX[7:0] = 8'b10010000;     // 9
  6'b001000: HEX[7:0] = 8'b10000000;     // 8
  6'b000111: HEX[7:0] = 8'b11111000;     // 7
  6'b000110: HEX[7:0] = 8'b10000010;     // 6
  6'b000101: HEX[7:0] = 8'b10010010;     // 5
  6'b000100: HEX[7:0] = 8'b10011001;     // 4
  6'b000011: HEX[7:0] = 8'b10110000;     // 3
  6'b000010: HEX[7:0] = 8'b10100100;     // 2
  6'b000001: HEX[7:0] = 8'b11111001;     // 1
  6'b000000: HEX[7:0] = 8'b11000000;     // 0  
  default: HEX[7:0] = 8'b11111111;
endcase 

endmodule