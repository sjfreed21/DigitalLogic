module top(ain, bin, cout);
    input ain, bin;
    output cout;
assign cout = ain & bin;

endmodule // topain, bin, cout);input ain, bin;